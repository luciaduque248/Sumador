library verilog;
use verilog.vl_types.all;
entity tablasum_vlg_vec_tst is
end tablasum_vlg_vec_tst;
