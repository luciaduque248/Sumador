library verilog;
use verilog.vl_types.all;
entity fulladder4Bits_vlg_vec_tst is
end fulladder4Bits_vlg_vec_tst;
