library verilog;
use verilog.vl_types.all;
entity testSumador_vlg_vec_tst is
end testSumador_vlg_vec_tst;
